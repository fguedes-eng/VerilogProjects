module VrDlatch_tb ();
reg D, G;
wire Q;


VrDlatch dut(D, G, Q);

initial begin
    

end

endmodule