module ShiftAdd_Multiplier (
    input clk,
    input rst,
    input [3:0] multiplier,
    input [3:0] multiplicand,
    input start,
    output [8:0] product,
    output done
);

    

endmodule